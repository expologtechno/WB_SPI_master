//List of Include Files

 `include "spi_base_test.sv"
 //`include "reset_test.sv"
 `include "lsb_8bit_data_test.sv"
 `include "ss_data_test.sv"
 `include "ie_data_test.sv"
 `include "miso_data_test.sv"
 `include "rand_data_test.sv"
