//`include "reset_seq.sv"
`include "sanity.sv"
`include "lsb_8bit_data.sv"
`include "miso_data.sv"
