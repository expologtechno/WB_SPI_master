//List of Include Files

 `include "spi_base_test.sv"
// `include "reset_test.sv"
 `include "lsb_8bit_data_test.sv"
 `include "lsb_16bit_data_test.sv"
 `include "lsb_32bit_data_test.sv"
 `include "lsb_64bit_data_test.sv"
 `include "lsb_128bit_data_test.sv"
 `include "msb_8bit_data_test.sv"
 `include "msb_16bit_data_test.sv"
 `include "msb_32bit_data_test.sv"
 `include "msb_64bit_data_test.sv"
 `include "msb_128bit_data_test.sv"
 `include "miso_data_test.sv"
 `include "Rx_raising_Tx_falling_test.sv"
 `include "Rx_falling_Tx_raising_test.sv"
