`include "reset_seq.sv"
`include "sanity.sv"
`include "lsb_8bit_data.sv"
`include "ss_data_seq.sv"
`include "ie_data_seq.sv"
`include "miso_data.sv"
`include "rand_data_seq.sv"
